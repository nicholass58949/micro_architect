// =============================================================================
// 文件名: output_buffer.v
// 功能: 输出数据缓存 - 存储计算结果
// 描述: 双端口RAM，支持激活函数单元写入和AXI读取
// =============================================================================

module output_buffer #(
    parameter DATA_WIDTH = 16,          // 数据位宽
    parameter BUFFER_DEPTH = 256,       // 缓存深度
    parameter ADDR_WIDTH = 8            // 地址位宽
)(
    // 时钟和复位
    input  wire                     clk,
    input  wire                     rst_n,
    
    // 写端口（来自激活函数单元）
    input  wire                     wr_en,
    input  wire [ADDR_WIDTH-1:0]    wr_addr,
    input  wire [DATA_WIDTH-1:0]    wr_data,
    
    // 读端口（到AXI接口）
    input  wire                     rd_en,
    input  wire [ADDR_WIDTH-1:0]    rd_addr,
    output reg  [DATA_WIDTH-1:0]    rd_data,
    output reg                      rd_valid
);

    // =========================================================================
    // 内部存储器
    // =========================================================================
    
    // 双端口RAM
    reg [DATA_WIDTH-1:0] buffer_mem [0:BUFFER_DEPTH-1];
    
    // 初始化
    integer i;
    initial begin
        for (i = 0; i < BUFFER_DEPTH; i = i + 1) begin
            buffer_mem[i] = {DATA_WIDTH{1'b0}};
        end
    end
    
    // =========================================================================
    // 写端口逻辑
    // =========================================================================
    
    always @(posedge clk) begin
        if (wr_en) begin
            buffer_mem[wr_addr] <= wr_data;
        end
    end
    
    // =========================================================================
    // 读端口逻辑
    // =========================================================================
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            rd_data <= {DATA_WIDTH{1'b0}};
            rd_valid <= 1'b0;
        end else begin
            if (rd_en) begin
                rd_data <= buffer_mem[rd_addr];
                rd_valid <= 1'b1;
            end else begin
                rd_valid <= 1'b0;
            end
        end
    end

endmodule

// =============================================================================
// 模块说明
// =============================================================================
//
// 功能描述：
// 输出缓存用于存储神经网络的计算结果（经过激活函数处理后的数据）。
// 采用双端口RAM设计，支持同时写入和读取操作。
//
// 工作原理：
// 1. 写端口：激活函数单元将处理后的数据写入缓存
// 2. 读端口：AXI接口从缓存读取结果返回给主机
// 3. 双端口设计允许写入和读取并行进行
//
// 存储容量：
// - 默认256个数据（可配置）
// - 每个数据16位（Q8.8格式）
// - 总容量：256 × 16 = 4096 bits = 512 bytes
//
// 接口协议：
// 写端口：
// - wr_en: 写使能，高电平有效
// - wr_addr: 写地址
// - wr_data: 写数据
//
// 读端口：
// - rd_en: 读使能，高电平有效
// - rd_addr: 读地址
// - rd_data: 读数据（下一周期有效）
// - rd_valid: 读数据有效标志
//
// 时序：
// - 写操作：同步写，数据在时钟上升沿写入
// - 读操作：同步读，数据在下一个时钟周期输出
// - 读延迟：1个时钟周期
//
// 数据流：
// 矩阵乘法单元 -> 激活函数单元 -> 输出缓存 -> AXI接口 -> 主机
//
// 使用场景：
// - 存储层输出结果
// - 中间层激活值（用于下一层计算）
// - 最终推理结果
//
// =============================================================================
