// =============================================================================
// 文件名: weight_buffer.v
// 功能: 权重缓存 - 存储神经网络权重数据
// 描述: 双端口RAM，支持AXI写入和矩阵乘法单元读取
// =============================================================================

module weight_buffer #(
    parameter DATA_WIDTH = 16,          // 数据位宽
    parameter BUFFER_DEPTH = 1024,      // 缓存深度（支持更大的权重矩阵）
    parameter ADDR_WIDTH = 10           // 地址位宽
)(
    // 时钟和复位
    input  wire                     clk,
    input  wire                     rst_n,
    
    // 写端口（来自AXI接口）
    input  wire                     wr_en,
    input  wire [ADDR_WIDTH-1:0]    wr_addr,
    input  wire [DATA_WIDTH-1:0]    wr_data,
    
    // 读端口（到矩阵乘法单元）
    input  wire                     rd_en,
    input  wire [ADDR_WIDTH-1:0]    rd_addr,
    output reg  [DATA_WIDTH-1:0]    rd_data,
    output reg                      rd_valid
);

    // =========================================================================
    // 内部存储器
    // =========================================================================
    
    // 双端口RAM
    reg [DATA_WIDTH-1:0] buffer_mem [0:BUFFER_DEPTH-1];
    
    // 初始化
    integer i;
    initial begin
        for (i = 0; i < BUFFER_DEPTH; i = i + 1) begin
            buffer_mem[i] = {DATA_WIDTH{1'b0}};
        end
    end
    
    // =========================================================================
    // 写端口逻辑
    // =========================================================================
    
    always @(posedge clk) begin
        if (wr_en) begin
            buffer_mem[wr_addr] <= wr_data;
        end
    end
    
    // =========================================================================
    // 读端口逻辑
    // =========================================================================
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            rd_data <= {DATA_WIDTH{1'b0}};
            rd_valid <= 1'b0;
        end else begin
            if (rd_en) begin
                rd_data <= buffer_mem[rd_addr];
                rd_valid <= 1'b1;
            end else begin
                rd_valid <= 1'b0;
            end
        end
    end

endmodule

// =============================================================================
// 模块说明
// =============================================================================
//
// 功能描述：
// 权重缓存用于存储神经网络的权重参数。
// 采用双端口RAM设计，支持同时写入和读取操作。
//
// 工作原理：
// 1. 写端口：AXI接口将权重数据写入缓存
// 2. 读端口：矩阵乘法单元从缓存读取权重进行计算
// 3. 权重数据通常在初始化时加载，计算过程中保持不变
//
// 存储容量：
// - 默认1024个数据（可配置）
// - 每个数据16位（Q8.8格式）
// - 总容量：1024 × 16 = 16384 bits = 2048 bytes
// - 可存储多个权重矩阵（如4个8×8矩阵）
//
// 接口协议：
// 写端口：
// - wr_en: 写使能，高电平有效
// - wr_addr: 写地址
// - wr_data: 写数据
//
// 读端口：
// - rd_en: 读使能，高电平有效
// - rd_addr: 读地址
// - rd_data: 读数据（下一周期有效）
// - rd_valid: 读数据有效标志
//
// 时序：
// - 写操作：同步写，数据在时钟上升沿写入
// - 读操作：同步读，数据在下一个时钟周期输出
// - 读延迟：1个时钟周期
//
// 权重组织：
// 对于8×8矩阵，权重按行优先顺序存储：
// - 地址0-7：第一行权重
// - 地址8-15：第二行权重
// - ...
// - 地址56-63：第八行权重
//
// 使用场景：
// - 存储全连接层权重
// - 存储卷积核参数
// - 多层网络权重缓存
//
// =============================================================================
