// =============================================================================
// 文件名: processing_element.v
// 功能: 处理单元（PE）- NPU的基本计算单元
// 描述: 执行乘累加（MAC）运算，是矩阵乘法的基本构建块
// =============================================================================

module processing_element #(
    parameter DATA_WIDTH = 16  // 数据位宽（Q8.8定点数格式）
)(
    // 时钟和复位
    input  wire                     clk,
    input  wire                     rst_n,
    
    // 控制信号
    input  wire                     enable,      // 使能信号
    input  wire                     clear_acc,   // 清除累加器
    
    // 数据输入
    input  wire [DATA_WIDTH-1:0]    data_in,     // 输入数据（激活值）
    input  wire [DATA_WIDTH-1:0]    weight_in,   // 权重数据
    
    // 数据输出
    output reg  [DATA_WIDTH-1:0]    data_out,    // 输出数据（传递给下一个PE）
    output reg  [2*DATA_WIDTH-1:0]  acc_out      // 累加结果输出
);

    // =========================================================================
    // 内部信号定义
    // =========================================================================
    
    // 乘法结果（扩展位宽以避免溢出）
    reg [2*DATA_WIDTH-1:0] mult_result;
    
    // 累加器（扩展位宽）
    reg [2*DATA_WIDTH-1:0] accumulator;
    
    // =========================================================================
    // 乘法运算
    // =========================================================================
    // 执行有符号乘法：data_in * weight_in
    // Q8.8 * Q8.8 = Q16.16（需要右移8位恢复到Q8.8格式）
    
    always @(*) begin
        mult_result = $signed(data_in) * $signed(weight_in);
    end
    
    // =========================================================================
    // 累加运算
    // =========================================================================
    // 累加器逻辑：实现 acc = acc + (data_in * weight_in)
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            accumulator <= {(2*DATA_WIDTH){1'b0}};
        end else if (clear_acc) begin
            // 清除累加器
            accumulator <= {(2*DATA_WIDTH){1'b0}};
        end else if (enable) begin
            // 累加新的乘法结果
            accumulator <= accumulator + mult_result;
        end
    end
    
    // =========================================================================
    // 数据流传递
    // =========================================================================
    // 将输入数据传递给下一个PE（用于脉动阵列）
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            data_out <= {DATA_WIDTH{1'b0}};
        end else if (enable) begin
            data_out <= data_in;
        end
    end
    
    // =========================================================================
    // 输出赋值
    // =========================================================================
    
    always @(posedge clk or negedge rst_n) begin
        if (!rst_n) begin
            acc_out <= {(2*DATA_WIDTH){1'b0}};
        end else begin
            acc_out <= accumulator;
        end
    end

endmodule

// =============================================================================
// 模块说明
// =============================================================================
// 
// 功能描述：
// 处理单元（PE）是NPU的基本计算单元，执行乘累加（MAC）运算。
// 多个PE可以组成脉动阵列，实现高效的矩阵乘法。
//
// 工作原理：
// 1. 接收输入数据（激活值）和权重数据
// 2. 执行乘法运算：mult_result = data_in * weight_in
// 3. 将乘法结果累加到累加器：accumulator += mult_result
// 4. 将输入数据传递给下一个PE（用于脉动阵列数据流）
//
// 数据格式：
// - 采用Q8.8定点数格式（8位整数 + 8位小数）
// - 乘法结果为Q16.16格式（需要后续处理）
// - 累加器使用32位宽度以避免溢出
//
// 时序：
// - 所有寄存器在时钟上升沿更新
// - 乘法运算为组合逻辑（当前周期完成）
// - 累加器在下一个时钟周期更新
//
// 控制信号：
// - enable: 高电平时PE工作，低电平时保持状态
// - clear_acc: 高电平时清除累加器，用于开始新的矩阵乘法
//
// 使用场景：
// - 矩阵乘法运算
// - 卷积运算
// - 全连接层计算
//
// =============================================================================
